`timescale 1ns / 1ps

module model_uart(/*AUTOARG*/
   // Outputs
   TX,
   // Inputs
   RX
   );

   output TX;
   input  RX;

   parameter baud    = 115200;
   parameter bittime = 1000000000/baud;
   parameter name    = "UART0";
   
   reg [7:0] rxData;
   reg [31:0] inputData;
   // have a bigger buffer to store any arbitrary amt of rx data, clear buffer by printing out when receive \r
   // 4 bytes, print out all 4 bytes when you see carriage return (2 bytes)
   event     evBit;
   event     evByte;
   event     evTxBit;
   event     evTxByte;
   reg       TX;

   initial
     begin
        TX = 1'b1;
     end
   
   always @ (negedge RX)
     begin
        rxData[7:0] = 8'h0;
        #(0.5*bittime);
        repeat (8)
          begin
             #bittime ->evBit;
             rxData[7:0] = {RX,rxData[7:1]};
          end
        ->evByte;
//        $display("%08x", rxData);
         if (rxData == 8'h0A)
            begin
               $display("%d %s Received word %08x (%c%c%c%c)", $stime, name,
                  inputData,
                  inputData[31:24],
                  inputData[23:16],
                  inputData[15:8],
                  inputData[7:0]);
               inputData[31:0] = 32'h0;
            end
         else
            begin
               inputData = {inputData[23:0], rxData};
            end
         // $display ("%d %s Received bytes %02x (%s)", $stime, name, rxData, rxData);
     end

   task tskRxData;
      output [7:0] data;
      begin
         @(evByte);
         data = rxData;
      end
   endtask // for
      
   task tskTxData;
      input [7:0] data;
      reg [9:0]   tmp;
      integer     i;
      begin
         tmp = {1'b1, data[7:0], 1'b0};
         for (i=0;i<10;i=i+1)
           begin
              TX = tmp[i];
              #bittime;
              ->evTxBit;
           end
         ->evTxByte;
      end
   endtask // tskTxData
   
endmodule // model_uart







